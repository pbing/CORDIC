/* arctan() for 17 iterations */
const bit signed [width + guard_bits - 3:0] atan_z[iterations] = '{65536, 38688, 20442, 10377, 5208, 2607, 1304, 652, 326, 163, 81, 41, 20, 10, 5, 3, 1};
