/* arctan() for 18 iterations */
const bit signed [width + guard_bits - 1:0] atan_z[iterations] = '{33'd1073741824, 33'd633866811, 33'd334917815, 33'd170009512, 33'd85334662, 33'd42708931, 33'd21359677, 33'd10680490, 33'd5340327, 33'd2670173, 33'd1335088, 33'd667544, 33'd333772, 33'd166886, 33'd83443, 33'd41722, 33'd20861, 33'd10430};
