/* arctan() for 18 iterations */
const bit signed [width + guard_bits - 1:0] atan_z[iterations] = '{262144, 154753, 81767, 41506, 20834, 10427, 5215, 2608, 1304, 652, 326, 163, 81, 41, 20, 10, 5, 3};
