/* arctan() for 19 iterations */
const bit signed [width + guard_bits - 1:0] atan_z[iterations] = '{35'd4294967296, 35'd2535467245, 35'd1339671259, 35'd680038049, 35'd341338648, 35'd170835723, 35'd85438707, 35'd42721961, 35'd21361306, 35'd10680694, 35'd5340352, 35'd2670177, 35'd1335088, 35'd667544, 35'd333772, 35'd166886, 35'd83443, 35'd41722, 35'd20861};
